module mongo

pub struct C.mongoc_client_t{}
pub struct C.mongoc_database_t{}
pub struct C.mongoc_collection_t{}
pub struct C.mongoc_uri_t{}