module mongo

#flag -I/usr/local/include/libmongoc-1.0
#flag -lmongoc-1.0
#include "mongoc/mongoc.h"

