module mongo

//
//	mongoc_*
//
struct C.mongoc_client_t{}
struct C.mongoc_database_t{}
struct C.mongoc_collection_t{}
struct C.mongoc_uri_t{}