module bson

#flag -I/usr/local/include/libbson-1.0
#flag -lbson-1.0
#include "bson/bson.h"
